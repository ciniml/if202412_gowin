tb_counter_8bit.sv